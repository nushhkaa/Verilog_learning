`timescale 1ns/1ns  
`include "test2.v"
//C:\iverilog\gtkwave\bin\gtkwave.exe
// module test2_tb;
// reg I;
// reg[1:0]S;
// wire [3:0]O;

// decoder_generate G1(O,I,S);
// initial begin
//     $display("First test started");
//     $monitor ($time, "    O = %b, I= %b, S = %h", O, I, S);
//     I = 1;      S = 0; #5
//     S = 1; #5
//     I = 0;      S = 0; #5
//     S = 1; #5
    
//     $display("First test complete");
//     $finish;
// end

// endmodule

module latchtest ;
reg 
    
endmodule